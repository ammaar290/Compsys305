LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.NUMERIC_STD.all;

ENTITY flappyBird IS
    PORT (
        pb1, pb2, clk, vert_sync : IN std_logic;
        pixel_row, pixel_column : IN std_logic_vector(9 DOWNTO 0);
        red, green, blue : OUT std_logic;
        collision_detected : OUT std_logic);
END flappyBird;

ARCHITECTURE behavior OF flappyBird IS
    -- Signals from Bird
    SIGNAL ball_on : std_logic;
    SIGNAL size : std_logic_vector(9 DOWNTO 0);  
    SIGNAL ball_y_pos : std_logic_vector(9 DOWNTO 0);
    SIGNAL ball_y_pos_T : std_logic_vector(9 DOWNTO 0);
    SIGNAL ball_x_pos : std_logic_vector(10 DOWNTO 0);
    SIGNAL ball_y_motion : std_logic_vector(9 DOWNTO 0);
    -- Signals from Pipes
    SIGNAL ball_on_upper, ball_on_lower : std_logic;
    SIGNAL sizex : std_logic_vector(9 DOWNTO 0);  
    SIGNAL ball_y_pos_upper, ball_y_pos_lower : std_logic_vector(9 DOWNTO 0);
    TYPE array_type is ARRAY (1 to 5) of std_logic_vector(9 DOWNTO 0);
    SIGNAL x_pos_arr : array_type;
    SIGNAL counter : integer range 0 to 333333 := 0;
    SIGNAL init_done: std_logic := '0';

BEGIN
    size <= std_logic_vector(to_unsigned(8,10));
    ball_x_pos <= std_logic_vector(to_unsigned(100,11));

 ball_on <= '1' when 
    (((unsigned('0' & ball_x_pos) <= (unsigned('0' & pixel_column) + unsigned(size))) and 
    (unsigned('0' & pixel_column) <= (unsigned('0' & ball_x_pos) + unsigned(size))) and 
    (unsigned('0' & ball_y_pos) <= (unsigned(pixel_row) + unsigned(size))) and 
    (unsigned('0' & pixel_row) <= (unsigned('0' & ball_y_pos) + unsigned(size)))
    else '0';

    Red <=  ball_on;
    Green <= ball_on;
    Blue <=  ball_on;

    sizex <= std_logic_vector(to_unsigned(20,10));  
    ball_y_pos_upper <= std_logic_vector(to_unsigned(150,10));
    ball_y_pos_lower <= std_logic_vector(to_unsigned(250,10));

    process (clk)
    begin
        if rising_edge(clk) then
            if init_done = '0' then
                x_pos_arr(1) <= std_logic_vector(to_unsigned(590,10));
                x_pos_arr(2) <= std_logic_vector(to_unsigned(480,10));
                x_pos_arr(3) <= std_logic_vector(to_unsigned(370,10));
                x_pos_arr(4) <= std_logic_vector(to_unsigned(260,10));
                x_pos_arr(5) <= std_logic_vector(to_unsigned(150,10));
                init_done <= '1';
            else
                counter <= counter + 1;
                if counter >= 333333 then
                    for i in 1 to 5 loop
                        if unsigned(x_pos_arr(i)) = 0 then
                            x_pos_arr(i) <= std_logic_vector(to_unsigned(800,10));
                        else
                            x_pos_arr(i) <= std_logic_vector(unsigned(x_pos_arr(i)) - 1);
                        end if;
                    end loop;
                    counter <= 0;
                end if;
            end if;
        end if;
    end process;

  process (pixel_row, pixel_column)
    begin
        ball_on_upper <= '0';
        ball_on_lower <= '0';
        for i in 1 to 5 loop
            if (( unsigned('0' & x_pos_arr(i)) <= unsigned(pixel_column))
                and (unsigned(pixel_column) < unsigned('0' & x_pos_arr(i)) + unsigned(sizex))) then
                if (unsigned(pixel_row) < unsigned(ball_y_pos_upper)) then
                    ball_on_upper <= '1';
                end if;
                if (unsigned(pixel_row) >= unsigned(ball_y_pos_lower)) then
                    ball_on_lower <= '1';
                end if;
            end if;
        end loop;
    end process;

    Move_Ball: process (vert_sync)  	
    begin
        if (rising_edge(vert_sync)) then
            if(pb1 = '1') then
                ball_y_motion <= std_logic_vector(to_unsigned(5,10));
            else
                ball_y_motion <= ball_y_motion - std_logic_vector(to_unsigned(1,10));
            end if;

            if(ball_y_pos <= "0111000010") then
                ball_y_pos_T <= "0110000000";
            else
                ball_y_pos_T <= ball_y_pos + ball_y_motion;
            end if;

            ball_y_pos <= ball_y_pos_T;
        end if;
    end process Move_Ball;

    collision_detected <= '1' when (ball_on = '1' and (ball_on_upper = '1' or ball_on_lower = '1')) else '0';

END behavior;
